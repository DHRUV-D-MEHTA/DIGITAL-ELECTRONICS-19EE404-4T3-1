library verilog;
use verilog.vl_types.all;
entity EX6_vlg_check_tst is
    port(
        q               : in     vl_logic;
        q_bar           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end EX6_vlg_check_tst;
