library verilog;
use verilog.vl_types.all;
entity EX5_vlg_vec_tst is
end EX5_vlg_vec_tst;
