library verilog;
use verilog.vl_types.all;
entity EX6_vlg_vec_tst is
end EX6_vlg_vec_tst;
