library verilog;
use verilog.vl_types.all;
entity EX5_vlg_check_tst is
    port(
        dout0           : in     vl_logic;
        dout1           : in     vl_logic;
        dout2           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end EX5_vlg_check_tst;
