library verilog;
use verilog.vl_types.all;
entity HALF_SUBTRACTOR_vlg_vec_tst is
end HALF_SUBTRACTOR_vlg_vec_tst;
