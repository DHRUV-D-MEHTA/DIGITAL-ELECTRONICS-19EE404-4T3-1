library verilog;
use verilog.vl_types.all;
entity HALF_ADDER_vlg_vec_tst is
end HALF_ADDER_vlg_vec_tst;
