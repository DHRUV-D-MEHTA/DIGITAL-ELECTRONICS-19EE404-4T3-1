library verilog;
use verilog.vl_types.all;
entity FULL_SUBTRACTOR_vlg_vec_tst is
end FULL_SUBTRACTOR_vlg_vec_tst;
