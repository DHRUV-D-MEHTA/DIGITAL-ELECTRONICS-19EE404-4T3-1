library verilog;
use verilog.vl_types.all;
entity EX11 is
    port(
        clk             : in     vl_logic;
        q1              : out    vl_logic;
        q2              : out    vl_logic;
        q3              : out    vl_logic
    );
end EX11;
