library verilog;
use verilog.vl_types.all;
entity EX10_vlg_check_tst is
    port(
        so              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end EX10_vlg_check_tst;
