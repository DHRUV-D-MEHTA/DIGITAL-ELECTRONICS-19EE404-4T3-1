library verilog;
use verilog.vl_types.all;
entity EX7_vlg_check_tst is
    port(
        q               : in     vl_logic;
        qb              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end EX7_vlg_check_tst;
