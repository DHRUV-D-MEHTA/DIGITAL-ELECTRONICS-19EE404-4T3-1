library verilog;
use verilog.vl_types.all;
entity EX8_vlg_vec_tst is
end EX8_vlg_vec_tst;
