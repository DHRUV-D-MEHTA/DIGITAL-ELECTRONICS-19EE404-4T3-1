library verilog;
use verilog.vl_types.all;
entity EX7_vlg_vec_tst is
end EX7_vlg_vec_tst;
