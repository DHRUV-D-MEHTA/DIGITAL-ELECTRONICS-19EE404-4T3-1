library verilog;
use verilog.vl_types.all;
entity EX5 is
    port(
        dout0           : out    vl_logic;
        dout1           : out    vl_logic;
        dout2           : out    vl_logic;
        din0            : in     vl_logic;
        din1            : in     vl_logic;
        din2            : in     vl_logic;
        din3            : in     vl_logic;
        din4            : in     vl_logic;
        din5            : in     vl_logic;
        din6            : in     vl_logic;
        din7            : in     vl_logic
    );
end EX5;
