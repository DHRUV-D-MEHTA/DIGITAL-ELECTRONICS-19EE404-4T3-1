library verilog;
use verilog.vl_types.all;
entity EX2_vlg_vec_tst is
end EX2_vlg_vec_tst;
