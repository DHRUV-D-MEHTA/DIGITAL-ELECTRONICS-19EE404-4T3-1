library verilog;
use verilog.vl_types.all;
entity EX11_vlg_vec_tst is
end EX11_vlg_vec_tst;
