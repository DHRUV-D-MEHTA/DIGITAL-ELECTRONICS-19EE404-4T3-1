library verilog;
use verilog.vl_types.all;
entity EX9_vlg_vec_tst is
end EX9_vlg_vec_tst;
