library verilog;
use verilog.vl_types.all;
entity EX12_vlg_vec_tst is
end EX12_vlg_vec_tst;
