library verilog;
use verilog.vl_types.all;
entity EX10_vlg_vec_tst is
end EX10_vlg_vec_tst;
