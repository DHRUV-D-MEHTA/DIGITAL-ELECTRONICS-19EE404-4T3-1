library verilog;
use verilog.vl_types.all;
entity EX1_vlg_vec_tst is
end EX1_vlg_vec_tst;
